.param W1=25u W2=29u W3=53u W4=32u W5=99u
.param W6=20u W7=15u